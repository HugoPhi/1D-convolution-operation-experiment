module top (
    
    );
    
endmodule
